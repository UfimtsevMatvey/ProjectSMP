//Myltiple steps adder add 128bit numbers
module two_step_adder64()

endmodule